module home_work3 (z, x, y);
output z;
input x;
input y;
assign z = x & y;
endmodule